`timescale 1ns / 1ps


module soc(

    );
endmodule
