`timescale 1ns / 1ps

`ifndef _DEFS_SV_
`define _DEFS_SV_

parameter WORD_SIZE = 32;
parameter ADDR_LEN = 5;


`endif